module tx(
    input clk,
    input n_rst,
    input 

);

